library verilog;
use verilog.vl_types.all;
entity ULAula_vlg_vec_tst is
end ULAula_vlg_vec_tst;
